magic
tech sky130A
magscale 1 2
timestamp 1659333009
<< obsli1 >>
rect 1104 2159 158884 157777
<< obsm1 >>
rect 14 2128 159146 157888
<< metal2 >>
rect 662 159200 718 160000
rect 7102 159200 7158 160000
rect 12898 159200 12954 160000
rect 18694 159200 18750 160000
rect 24490 159200 24546 160000
rect 30286 159200 30342 160000
rect 36082 159200 36138 160000
rect 41878 159200 41934 160000
rect 48318 159200 48374 160000
rect 54114 159200 54170 160000
rect 59910 159200 59966 160000
rect 65706 159200 65762 160000
rect 71502 159200 71558 160000
rect 77298 159200 77354 160000
rect 83738 159200 83794 160000
rect 89534 159200 89590 160000
rect 95330 159200 95386 160000
rect 101126 159200 101182 160000
rect 106922 159200 106978 160000
rect 112718 159200 112774 160000
rect 118514 159200 118570 160000
rect 124954 159200 125010 160000
rect 130750 159200 130806 160000
rect 136546 159200 136602 160000
rect 142342 159200 142398 160000
rect 148138 159200 148194 160000
rect 153934 159200 153990 160000
rect 159730 159200 159786 160000
rect 18 0 74 800
rect 5814 0 5870 800
rect 11610 0 11666 800
rect 17406 0 17462 800
rect 23202 0 23258 800
rect 28998 0 29054 800
rect 34794 0 34850 800
rect 41234 0 41290 800
rect 47030 0 47086 800
rect 52826 0 52882 800
rect 58622 0 58678 800
rect 64418 0 64474 800
rect 70214 0 70270 800
rect 76010 0 76066 800
rect 82450 0 82506 800
rect 88246 0 88302 800
rect 94042 0 94098 800
rect 99838 0 99894 800
rect 105634 0 105690 800
rect 111430 0 111486 800
rect 117870 0 117926 800
rect 123666 0 123722 800
rect 129462 0 129518 800
rect 135258 0 135314 800
rect 141054 0 141110 800
rect 146850 0 146906 800
rect 152646 0 152702 800
rect 159086 0 159142 800
<< obsm2 >>
rect 20 159144 606 159338
rect 774 159144 7046 159338
rect 7214 159144 12842 159338
rect 13010 159144 18638 159338
rect 18806 159144 24434 159338
rect 24602 159144 30230 159338
rect 30398 159144 36026 159338
rect 36194 159144 41822 159338
rect 41990 159144 48262 159338
rect 48430 159144 54058 159338
rect 54226 159144 59854 159338
rect 60022 159144 65650 159338
rect 65818 159144 71446 159338
rect 71614 159144 77242 159338
rect 77410 159144 83682 159338
rect 83850 159144 89478 159338
rect 89646 159144 95274 159338
rect 95442 159144 101070 159338
rect 101238 159144 106866 159338
rect 107034 159144 112662 159338
rect 112830 159144 118458 159338
rect 118626 159144 124898 159338
rect 125066 159144 130694 159338
rect 130862 159144 136490 159338
rect 136658 159144 142286 159338
rect 142454 159144 148082 159338
rect 148250 159144 153878 159338
rect 154046 159144 159140 159338
rect 20 856 159140 159144
rect 130 800 5758 856
rect 5926 800 11554 856
rect 11722 800 17350 856
rect 17518 800 23146 856
rect 23314 800 28942 856
rect 29110 800 34738 856
rect 34906 800 41178 856
rect 41346 800 46974 856
rect 47142 800 52770 856
rect 52938 800 58566 856
rect 58734 800 64362 856
rect 64530 800 70158 856
rect 70326 800 75954 856
rect 76122 800 82394 856
rect 82562 800 88190 856
rect 88358 800 93986 856
rect 94154 800 99782 856
rect 99950 800 105578 856
rect 105746 800 111374 856
rect 111542 800 117814 856
rect 117982 800 123610 856
rect 123778 800 129406 856
rect 129574 800 135202 856
rect 135370 800 140998 856
rect 141166 800 146794 856
rect 146962 800 152590 856
rect 152758 800 159030 856
<< metal3 >>
rect 0 155048 800 155168
rect 159200 153688 160000 153808
rect 0 148928 800 149048
rect 159200 147568 160000 147688
rect 0 142808 800 142928
rect 159200 141448 160000 141568
rect 0 136688 800 136808
rect 159200 135328 160000 135448
rect 0 130568 800 130688
rect 159200 129208 160000 129328
rect 0 124448 800 124568
rect 159200 123088 160000 123208
rect 0 117648 800 117768
rect 159200 116288 160000 116408
rect 0 111528 800 111648
rect 159200 110168 160000 110288
rect 0 105408 800 105528
rect 159200 104048 160000 104168
rect 0 99288 800 99408
rect 159200 97928 160000 98048
rect 0 93168 800 93288
rect 159200 91808 160000 91928
rect 0 87048 800 87168
rect 159200 85688 160000 85808
rect 0 80248 800 80368
rect 159200 79568 160000 79688
rect 0 74128 800 74248
rect 159200 72768 160000 72888
rect 0 68008 800 68128
rect 159200 66648 160000 66768
rect 0 61888 800 62008
rect 159200 60528 160000 60648
rect 0 55768 800 55888
rect 159200 54408 160000 54528
rect 0 49648 800 49768
rect 159200 48288 160000 48408
rect 0 43528 800 43648
rect 159200 42168 160000 42288
rect 0 36728 800 36848
rect 159200 35368 160000 35488
rect 0 30608 800 30728
rect 159200 29248 160000 29368
rect 0 24488 800 24608
rect 159200 23128 160000 23248
rect 0 18368 800 18488
rect 159200 17008 160000 17128
rect 0 12248 800 12368
rect 159200 10888 160000 11008
rect 0 6128 800 6248
rect 159200 4768 160000 4888
<< obsm3 >>
rect 800 155248 159200 157793
rect 880 154968 159200 155248
rect 800 153888 159200 154968
rect 800 153608 159120 153888
rect 800 149128 159200 153608
rect 880 148848 159200 149128
rect 800 147768 159200 148848
rect 800 147488 159120 147768
rect 800 143008 159200 147488
rect 880 142728 159200 143008
rect 800 141648 159200 142728
rect 800 141368 159120 141648
rect 800 136888 159200 141368
rect 880 136608 159200 136888
rect 800 135528 159200 136608
rect 800 135248 159120 135528
rect 800 130768 159200 135248
rect 880 130488 159200 130768
rect 800 129408 159200 130488
rect 800 129128 159120 129408
rect 800 124648 159200 129128
rect 880 124368 159200 124648
rect 800 123288 159200 124368
rect 800 123008 159120 123288
rect 800 117848 159200 123008
rect 880 117568 159200 117848
rect 800 116488 159200 117568
rect 800 116208 159120 116488
rect 800 111728 159200 116208
rect 880 111448 159200 111728
rect 800 110368 159200 111448
rect 800 110088 159120 110368
rect 800 105608 159200 110088
rect 880 105328 159200 105608
rect 800 104248 159200 105328
rect 800 103968 159120 104248
rect 800 99488 159200 103968
rect 880 99208 159200 99488
rect 800 98128 159200 99208
rect 800 97848 159120 98128
rect 800 93368 159200 97848
rect 880 93088 159200 93368
rect 800 92008 159200 93088
rect 800 91728 159120 92008
rect 800 87248 159200 91728
rect 880 86968 159200 87248
rect 800 85888 159200 86968
rect 800 85608 159120 85888
rect 800 80448 159200 85608
rect 880 80168 159200 80448
rect 800 79768 159200 80168
rect 800 79488 159120 79768
rect 800 74328 159200 79488
rect 880 74048 159200 74328
rect 800 72968 159200 74048
rect 800 72688 159120 72968
rect 800 68208 159200 72688
rect 880 67928 159200 68208
rect 800 66848 159200 67928
rect 800 66568 159120 66848
rect 800 62088 159200 66568
rect 880 61808 159200 62088
rect 800 60728 159200 61808
rect 800 60448 159120 60728
rect 800 55968 159200 60448
rect 880 55688 159200 55968
rect 800 54608 159200 55688
rect 800 54328 159120 54608
rect 800 49848 159200 54328
rect 880 49568 159200 49848
rect 800 48488 159200 49568
rect 800 48208 159120 48488
rect 800 43728 159200 48208
rect 880 43448 159200 43728
rect 800 42368 159200 43448
rect 800 42088 159120 42368
rect 800 36928 159200 42088
rect 880 36648 159200 36928
rect 800 35568 159200 36648
rect 800 35288 159120 35568
rect 800 30808 159200 35288
rect 880 30528 159200 30808
rect 800 29448 159200 30528
rect 800 29168 159120 29448
rect 800 24688 159200 29168
rect 880 24408 159200 24688
rect 800 23328 159200 24408
rect 800 23048 159120 23328
rect 800 18568 159200 23048
rect 880 18288 159200 18568
rect 800 17208 159200 18288
rect 800 16928 159120 17208
rect 800 12448 159200 16928
rect 880 12168 159200 12448
rect 800 11088 159200 12168
rect 800 10808 159120 11088
rect 800 6328 159200 10808
rect 880 6048 159200 6328
rect 800 4968 159200 6048
rect 800 4688 159120 4968
rect 800 2143 159200 4688
<< metal4 >>
rect 4208 2128 4528 157808
rect 19568 2128 19888 157808
rect 34928 2128 35248 157808
rect 50288 2128 50608 157808
rect 65648 2128 65968 157808
rect 81008 2128 81328 157808
rect 96368 2128 96688 157808
rect 111728 2128 112048 157808
rect 127088 2128 127408 157808
rect 142448 2128 142768 157808
rect 157808 2128 158128 157808
<< obsm4 >>
rect 20299 8875 34848 157589
rect 35328 8875 50208 157589
rect 50688 8875 65568 157589
rect 66048 8875 80928 157589
rect 81408 8875 96288 157589
rect 96768 8875 111648 157589
rect 112128 8875 127008 157589
rect 127488 8875 133893 157589
<< labels >>
rlabel metal2 s 18694 159200 18750 160000 6 clock
port 1 nsew signal input
rlabel metal2 s 141054 0 141110 800 6 io_wbs_ack_o
port 2 nsew signal output
rlabel metal3 s 159200 129208 160000 129328 6 io_wbs_adr_i[0]
port 3 nsew signal input
rlabel metal3 s 0 93168 800 93288 6 io_wbs_adr_i[10]
port 4 nsew signal input
rlabel metal3 s 0 105408 800 105528 6 io_wbs_adr_i[11]
port 5 nsew signal input
rlabel metal2 s 101126 159200 101182 160000 6 io_wbs_adr_i[12]
port 6 nsew signal input
rlabel metal2 s 118514 159200 118570 160000 6 io_wbs_adr_i[13]
port 7 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 io_wbs_adr_i[14]
port 8 nsew signal input
rlabel metal3 s 0 74128 800 74248 6 io_wbs_adr_i[15]
port 9 nsew signal input
rlabel metal3 s 159200 110168 160000 110288 6 io_wbs_adr_i[16]
port 10 nsew signal input
rlabel metal3 s 159200 85688 160000 85808 6 io_wbs_adr_i[17]
port 11 nsew signal input
rlabel metal3 s 159200 4768 160000 4888 6 io_wbs_adr_i[18]
port 12 nsew signal input
rlabel metal3 s 0 124448 800 124568 6 io_wbs_adr_i[19]
port 13 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 io_wbs_adr_i[1]
port 14 nsew signal input
rlabel metal2 s 135258 0 135314 800 6 io_wbs_adr_i[20]
port 15 nsew signal input
rlabel metal3 s 159200 35368 160000 35488 6 io_wbs_adr_i[21]
port 16 nsew signal input
rlabel metal2 s 83738 159200 83794 160000 6 io_wbs_adr_i[22]
port 17 nsew signal input
rlabel metal3 s 0 136688 800 136808 6 io_wbs_adr_i[23]
port 18 nsew signal input
rlabel metal2 s 48318 159200 48374 160000 6 io_wbs_adr_i[24]
port 19 nsew signal input
rlabel metal3 s 159200 147568 160000 147688 6 io_wbs_adr_i[25]
port 20 nsew signal input
rlabel metal2 s 95330 159200 95386 160000 6 io_wbs_adr_i[26]
port 21 nsew signal input
rlabel metal3 s 159200 29248 160000 29368 6 io_wbs_adr_i[27]
port 22 nsew signal input
rlabel metal3 s 0 87048 800 87168 6 io_wbs_adr_i[28]
port 23 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 io_wbs_adr_i[29]
port 24 nsew signal input
rlabel metal3 s 0 55768 800 55888 6 io_wbs_adr_i[2]
port 25 nsew signal input
rlabel metal3 s 159200 23128 160000 23248 6 io_wbs_adr_i[30]
port 26 nsew signal input
rlabel metal2 s 112718 159200 112774 160000 6 io_wbs_adr_i[31]
port 27 nsew signal input
rlabel metal3 s 0 111528 800 111648 6 io_wbs_adr_i[3]
port 28 nsew signal input
rlabel metal2 s 34794 0 34850 800 6 io_wbs_adr_i[4]
port 29 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 io_wbs_adr_i[5]
port 30 nsew signal input
rlabel metal2 s 148138 159200 148194 160000 6 io_wbs_adr_i[6]
port 31 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 io_wbs_adr_i[7]
port 32 nsew signal input
rlabel metal3 s 0 30608 800 30728 6 io_wbs_adr_i[8]
port 33 nsew signal input
rlabel metal2 s 159730 159200 159786 160000 6 io_wbs_adr_i[9]
port 34 nsew signal input
rlabel metal2 s 130750 159200 130806 160000 6 io_wbs_cyc_i
port 35 nsew signal input
rlabel metal3 s 159200 135328 160000 135448 6 io_wbs_dat_i[0]
port 36 nsew signal input
rlabel metal3 s 159200 153688 160000 153808 6 io_wbs_dat_i[10]
port 37 nsew signal input
rlabel metal3 s 159200 66648 160000 66768 6 io_wbs_dat_i[11]
port 38 nsew signal input
rlabel metal3 s 159200 54408 160000 54528 6 io_wbs_dat_i[12]
port 39 nsew signal input
rlabel metal2 s 54114 159200 54170 160000 6 io_wbs_dat_i[13]
port 40 nsew signal input
rlabel metal2 s 59910 159200 59966 160000 6 io_wbs_dat_i[14]
port 41 nsew signal input
rlabel metal3 s 159200 123088 160000 123208 6 io_wbs_dat_i[15]
port 42 nsew signal input
rlabel metal2 s 77298 159200 77354 160000 6 io_wbs_dat_i[16]
port 43 nsew signal input
rlabel metal2 s 41234 0 41290 800 6 io_wbs_dat_i[17]
port 44 nsew signal input
rlabel metal2 s 65706 159200 65762 160000 6 io_wbs_dat_i[18]
port 45 nsew signal input
rlabel metal2 s 159086 0 159142 800 6 io_wbs_dat_i[19]
port 46 nsew signal input
rlabel metal2 s 89534 159200 89590 160000 6 io_wbs_dat_i[1]
port 47 nsew signal input
rlabel metal3 s 0 117648 800 117768 6 io_wbs_dat_i[20]
port 48 nsew signal input
rlabel metal2 s 41878 159200 41934 160000 6 io_wbs_dat_i[21]
port 49 nsew signal input
rlabel metal3 s 159200 10888 160000 11008 6 io_wbs_dat_i[22]
port 50 nsew signal input
rlabel metal3 s 159200 141448 160000 141568 6 io_wbs_dat_i[23]
port 51 nsew signal input
rlabel metal2 s 136546 159200 136602 160000 6 io_wbs_dat_i[24]
port 52 nsew signal input
rlabel metal2 s 117870 0 117926 800 6 io_wbs_dat_i[25]
port 53 nsew signal input
rlabel metal2 s 58622 0 58678 800 6 io_wbs_dat_i[26]
port 54 nsew signal input
rlabel metal3 s 159200 42168 160000 42288 6 io_wbs_dat_i[27]
port 55 nsew signal input
rlabel metal3 s 0 61888 800 62008 6 io_wbs_dat_i[28]
port 56 nsew signal input
rlabel metal3 s 0 80248 800 80368 6 io_wbs_dat_i[29]
port 57 nsew signal input
rlabel metal2 s 152646 0 152702 800 6 io_wbs_dat_i[2]
port 58 nsew signal input
rlabel metal2 s 30286 159200 30342 160000 6 io_wbs_dat_i[30]
port 59 nsew signal input
rlabel metal2 s 123666 0 123722 800 6 io_wbs_dat_i[31]
port 60 nsew signal input
rlabel metal3 s 0 148928 800 149048 6 io_wbs_dat_i[3]
port 61 nsew signal input
rlabel metal3 s 0 24488 800 24608 6 io_wbs_dat_i[4]
port 62 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 io_wbs_dat_i[5]
port 63 nsew signal input
rlabel metal2 s 47030 0 47086 800 6 io_wbs_dat_i[6]
port 64 nsew signal input
rlabel metal2 s 146850 0 146906 800 6 io_wbs_dat_i[7]
port 65 nsew signal input
rlabel metal3 s 159200 79568 160000 79688 6 io_wbs_dat_i[8]
port 66 nsew signal input
rlabel metal3 s 159200 48288 160000 48408 6 io_wbs_dat_i[9]
port 67 nsew signal input
rlabel metal2 s 111430 0 111486 800 6 io_wbs_dat_o[0]
port 68 nsew signal output
rlabel metal3 s 0 130568 800 130688 6 io_wbs_dat_o[10]
port 69 nsew signal output
rlabel metal3 s 0 99288 800 99408 6 io_wbs_dat_o[11]
port 70 nsew signal output
rlabel metal3 s 0 36728 800 36848 6 io_wbs_dat_o[12]
port 71 nsew signal output
rlabel metal3 s 159200 60528 160000 60648 6 io_wbs_dat_o[13]
port 72 nsew signal output
rlabel metal3 s 159200 104048 160000 104168 6 io_wbs_dat_o[14]
port 73 nsew signal output
rlabel metal2 s 129462 0 129518 800 6 io_wbs_dat_o[15]
port 74 nsew signal output
rlabel metal3 s 159200 116288 160000 116408 6 io_wbs_dat_o[16]
port 75 nsew signal output
rlabel metal2 s 76010 0 76066 800 6 io_wbs_dat_o[17]
port 76 nsew signal output
rlabel metal2 s 662 159200 718 160000 6 io_wbs_dat_o[18]
port 77 nsew signal output
rlabel metal3 s 0 68008 800 68128 6 io_wbs_dat_o[19]
port 78 nsew signal output
rlabel metal2 s 18 0 74 800 6 io_wbs_dat_o[1]
port 79 nsew signal output
rlabel metal2 s 94042 0 94098 800 6 io_wbs_dat_o[20]
port 80 nsew signal output
rlabel metal2 s 24490 159200 24546 160000 6 io_wbs_dat_o[21]
port 81 nsew signal output
rlabel metal2 s 71502 159200 71558 160000 6 io_wbs_dat_o[22]
port 82 nsew signal output
rlabel metal3 s 0 18368 800 18488 6 io_wbs_dat_o[23]
port 83 nsew signal output
rlabel metal3 s 0 155048 800 155168 6 io_wbs_dat_o[24]
port 84 nsew signal output
rlabel metal2 s 23202 0 23258 800 6 io_wbs_dat_o[25]
port 85 nsew signal output
rlabel metal2 s 5814 0 5870 800 6 io_wbs_dat_o[26]
port 86 nsew signal output
rlabel metal2 s 142342 159200 142398 160000 6 io_wbs_dat_o[27]
port 87 nsew signal output
rlabel metal2 s 106922 159200 106978 160000 6 io_wbs_dat_o[28]
port 88 nsew signal output
rlabel metal2 s 70214 0 70270 800 6 io_wbs_dat_o[29]
port 89 nsew signal output
rlabel metal2 s 153934 159200 153990 160000 6 io_wbs_dat_o[2]
port 90 nsew signal output
rlabel metal3 s 159200 17008 160000 17128 6 io_wbs_dat_o[30]
port 91 nsew signal output
rlabel metal2 s 7102 159200 7158 160000 6 io_wbs_dat_o[31]
port 92 nsew signal output
rlabel metal3 s 159200 91808 160000 91928 6 io_wbs_dat_o[3]
port 93 nsew signal output
rlabel metal2 s 28998 0 29054 800 6 io_wbs_dat_o[4]
port 94 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 io_wbs_dat_o[5]
port 95 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 io_wbs_dat_o[6]
port 96 nsew signal output
rlabel metal3 s 159200 97928 160000 98048 6 io_wbs_dat_o[7]
port 97 nsew signal output
rlabel metal2 s 88246 0 88302 800 6 io_wbs_dat_o[8]
port 98 nsew signal output
rlabel metal3 s 0 43528 800 43648 6 io_wbs_dat_o[9]
port 99 nsew signal output
rlabel metal2 s 124954 159200 125010 160000 6 io_wbs_sel_i[0]
port 100 nsew signal input
rlabel metal2 s 12898 159200 12954 160000 6 io_wbs_sel_i[1]
port 101 nsew signal input
rlabel metal2 s 36082 159200 36138 160000 6 io_wbs_sel_i[2]
port 102 nsew signal input
rlabel metal2 s 105634 0 105690 800 6 io_wbs_sel_i[3]
port 103 nsew signal input
rlabel metal3 s 0 49648 800 49768 6 io_wbs_stb_i
port 104 nsew signal input
rlabel metal3 s 0 142808 800 142928 6 io_wbs_we_i
port 105 nsew signal input
rlabel metal3 s 159200 72768 160000 72888 6 reset
port 106 nsew signal input
rlabel metal4 s 4208 2128 4528 157808 6 vccd1
port 107 nsew power input
rlabel metal4 s 34928 2128 35248 157808 6 vccd1
port 107 nsew power input
rlabel metal4 s 65648 2128 65968 157808 6 vccd1
port 107 nsew power input
rlabel metal4 s 96368 2128 96688 157808 6 vccd1
port 107 nsew power input
rlabel metal4 s 127088 2128 127408 157808 6 vccd1
port 107 nsew power input
rlabel metal4 s 157808 2128 158128 157808 6 vccd1
port 107 nsew power input
rlabel metal4 s 19568 2128 19888 157808 6 vssd1
port 108 nsew ground input
rlabel metal4 s 50288 2128 50608 157808 6 vssd1
port 108 nsew ground input
rlabel metal4 s 81008 2128 81328 157808 6 vssd1
port 108 nsew ground input
rlabel metal4 s 111728 2128 112048 157808 6 vssd1
port 108 nsew ground input
rlabel metal4 s 142448 2128 142768 157808 6 vssd1
port 108 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 160000 160000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 34986764
string GDS_FILE /home/faiek/caravel_AES/caravel_AES/openlane/aes/runs/aes/results/finishing/aes.magic.gds
string GDS_START 1167592
<< end >>

